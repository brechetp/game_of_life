-- cellular automata.
-- computes the generation g+1 from the generation g on a window
--                WIDTH
-- ------------------------------------------------
-- |      N_CELL                                  |
-- |     --------                                 | HEIGHT
-- |     |      | 3 rows                          |
-- |     --------                                 |
-- |        |                                     |
-- |        v                                     |
-- ------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library celloux_lib;
use celloux_lib.pack_cell.all;
library WORK;
use WORK.main_pkg.all;

entity cell_ctrl is
  port(
    clk, rstn: in std_ulogic; -- clock and synchronous reset
    -- read / write signals to start reading / writing
    DONE_READING:  in std_ulogic; -- read_cell_vector is ready to be read
    DONE_WRITING: in std_ulogic; -- write_cell_vector is ready to be written, it has been written into mem
    READY_READING: out std_ulogic; -- the read_cell_vector has been read, it can now be changed by ADDR_CTR
    READY_WRITING: out std_ulogic; -- the write_cell_vector is ready to be written in memory
    -- n state of the world, 3 rows at a time of width BUFFER_SIZE
    read_cell_vector: in CELL_VECTOR(0 to N_CELL-1); -- read cells from memory
                                                                -- we only need this one as our window is gliding

    -- n+1 state of the world to be written in memory
    write_cell_vector:     out CELL_VECTOR(0 to N_CELL-3) -- cells to be written to memory
                                      -- this is the north register
    -- lock: out std_ulogic
  );
end entity cell_ctrl;

architecture arc of cell_ctrl is

  signal cells: window; -- the cells translated from the colors, 3 x N_CELL
  signal new_cells: CELL_VECTOR(0 to N_CELL-1);
  --signal -- new_data: std_logic := 'L';
  signal state: CELL_CTRL_STATE := FREEZE;

begin

  -- lock <= new_data;

  state_process: process(clk)
  begin
    if clk = '1' then
      if rstn = '0' then
        state <= FREEZE;
      else
        case state is
          when FREEZE =>
            if DONE_WRITING = '1' and DONE_READING = '1' then
              state <= NORMAL;
            else
              if DONE_WRITING = '1' then
                state <= WRITE;
              else
                if DONE_READING = '1' then
                  state <= READ;
                end if;
              end if;
            end if;

          when READ =>
            if DONE_READING = '0' then
              if DONE_WRITING = '1' then
                state <= WRITE;
              else
                state <= FREEZE;
              end if;
            else -- DONE_READING = '0'
              if DONE_WRITING = '1' then
                state <= NORMAL;
              end if;
            end if;

          when WRITE =>
            if DONE_WRITING = '0' then
              if DONE_READING = '1' then
                state <= READ;
              else
                state <= FREEZE;
              end if;
            else
              if DONE_READING = '1' then
                state <= NORMAL;
              end if;
            end if;

          when NORMAL => 
            if done_writing = '0' then
              if done_reading = '0' then
                state <= FREEZE;
              else
                state <= READ;
              end if;
            else
              if done_reading = '0' then
                state <= WRITE;
              end if;
            end if;
        end case;
      end if;
    end if;
  end process state_process;

            

  
  input: process(clk)
  begin
    if clk = '1' then
      if rstn = '0' then
        for i in 0 to N_CELL-1 loop
          cells(0, i) <= DEAD;
          cells(1, i) <= DEAD;
          cells(2, i) <= DEAD;
        end loop;
        READY_READING <= '0';
        -- new_data <= 'L';
      else
        READY_READING <= '0'; -- unless we say so, the memory is not ready to be overwritten
        if (state = READ) or (state = NORMAL) then -- we can't do anything unless the past generation has been written to memory
          for i in 0 to ( N_CELL-1 ) loop -- we slide the widow towards the south
            cells(0,i) <= cells(1,i);
            cells(1,i) <= cells(2,i);
            cells(2,i)  <= (read_cell_vector(i));
          end loop;
          READY_READING <= '1'; -- tells the mem the read_cell_vector has been read (it can be written), DONE_READING will be set to 0
          -- new_data <= 'H'; -- we can trust the computation of the generation g
        end if;
      end if; -- end of the reset block
    end if; -- end of the synchronous block
  end process input;


  GEN: for i in 1 to ( N_CELL-2 ) generate -- we create N_CELL-2 cells, mapped with each others
    CELL: entity CELLOUX_LIB.CELL(syn)
    port map(clk, rstn, '1', cells(0,i), cells(0,i+1), cells(1,i+1), cells(2,i+1), cells(2,i), cells(2,i-1), cells(1,i-1), cells(0,i-1), cells(1, i), new_cells(i));
  end generate GEN;

  output: process(clk)
  begin
    if clk = '1' then
      if rstn = '0' then
        for i in 0 to N_CELL-3 loop
          write_cell_vector(i) <= DEAD;
        end loop;
        READY_WRITING <= '0';
      else
        READY_WRITING <= '0'; -- we set READY_WRITING to 0 unless we cache the new cells in the write_cell_vector
        if (state = WRITE or state = NORMAL) then -- checks if new data is to be output and if the old one has been written
          for i in 0 to ( N_CELL-3 ) loop
            write_cell_vector(i) <= new_cells(i); -- output the soon-to-be-written cells
          end loop;
          READY_WRITING <= '1'; -- the DONE_WRITING will be set to 0 by address controller ?
          -- new_data <= 'L'; -- resolved type
        end if;
      end if; -- end of the reset block
    end if;-- end of the syncronous block
  end process;

end;

